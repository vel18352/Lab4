module tabla_6(input wire A,B,C, output wire Y);

  assign Y = ~B | C;
              
endmodule


