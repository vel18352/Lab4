module tabla_2(input wire A,B,C, output wire Y);

  assign Y = ~B;
              
endmodule


